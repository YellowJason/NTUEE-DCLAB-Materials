module Keyboard(
    input i_clk,
    input i_rst_n,
    // PS2 input signal
    input i_data,
    input i_ps2_clk,
    
    output [3:0] o_num1,
    output [3:0] o_num2
);


endmodule

module altpll (
	clk_clk,
	reset_reset_n,
	altpll_25_clk,
	altpll_65_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		altpll_25_clk;
	output		altpll_65_clk;
endmodule
